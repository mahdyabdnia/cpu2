module control(ins,reg2loc,uncondbr,br,MemRead,MemToReg,ALUOp,MemWrite,ALUsrc,RegWrite)
input reg2loc;



endmodule
