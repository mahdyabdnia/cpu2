module finaltestbench;
clock clk();
testbench2 tb2();

endmodule
